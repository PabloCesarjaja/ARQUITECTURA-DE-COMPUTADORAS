// Definir modulo y sus entradas y salidas
module _and (input A, input B, output C);//guion bajo mayusculas o minusculas
//2. declara señales/elementos internos
//NA
//3. comportamiento del modulo (asignaciones, instancias, conexiones)
assign C = A&B;



endmodule